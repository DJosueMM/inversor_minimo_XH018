*nmos minimo.sp

.subckt nmos g d

xm0 d g gnd! gnd! ne w=360n l=180n as=1.728e-13 ad=1.728e-13 ps=1.68e-06 pd=1.68e-06
+ nrs=0.75 nrd=0.75 m='1*1' par1='1*1' xf_subext=0

.ends
